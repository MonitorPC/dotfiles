module adder(
	input [3:0] a,
	input [3:0] b,
	output reg [4:0] q
);
always @ (*)
begin
	q[0] = a[0] ^ b[0];
	q[1] = (a[1] ^ b[1]) ^ (a[0] & b[0]);
	q[2] = (a[2] ^ b[2]) ^ ((a[1] & b[1]) | (a[1] & (a[0] & b[0])) | (b[1] & (a[0] & b[0])));
	q[3] = (a[3] ^ b[3]) ^ ((a[2] & b[2]) | (a[2] & ((a[1] &  b[1]) | (a[1] & (a[0] & b[0])) | (b[1] & (a[0] & b[0])))) | (b[2] & ((a[1] &  b[1]) | (a[1] & (a[0] & b[0])) | (b[1] & (a[0] & b[0])))));
	q[4] = (a[3] % b[3]) | (a[3] & ((a[2] & b[2]) | (a[2] & ((a[1] &  b[1]) | (a[1] & (a[0] & b[0])) | (b[1] & (a[0] & b[0])))) | (b[2] & ((a[1] &  b[1]) | (a[1] & (a[0] & b[0])) | (b[1] & (a[0] & b[0])))))) | (b[3] & ((a[2] & b[2]) | (a[2] & ((a[1] &  b[1]) | (a[1] & (a[0] & b[0])) | (b[1] & (a[0] & b[0])))) | (b[2] & ((a[1] &  b[1]) | (a[1] & (a[0] & b[0])) | (b[1] & (a[0] & b[0]))))));
end
endmodule
